netcdf drydep_tables {
dimensions:
  n_species_table = 131;
  NHen  = 6;
  chars = 16;
variables:
  
  char species_name_table(n_species_table,chars);
    species_name_table:long_name = "names of species in dry deposition tables" ;
  double dfoxd(n_species_table);
    dfoxd:long_name = "data for foxd (reactivity factor for oxidation)";
  double dheff(n_species_table,NHen);
    dheff:long_name = "data for effective Henry's Law coefficient";
  double mol_wghts(n_species_table);
    mol_wghts:long_name = "species molecular mass";
    mol_wghts:units = "grams/mole";
    
// global attributes:

  :Created_by = "Elizabeth Lundgren (Harvard University)";
  :Source = "GEOS-Chem version 14.3. gas-phase dry deposited species";

data:

  species_name_table =
         "ACET            ",
         "ACTA            ",
         "ALD2            ",
         "AROMP4          ",
         "AROMP5          ",
         "ATOOH           ",
         "BALD            ",
         "BENZP           ",
         "BR2             ",
         "BRCL            ",
         "BRNO3           ",
         "BZCO3H          ",
         "BZPAN           ",
         "CH2O            ",
         "CL2             ",
         "CLNO2           ",
         "CLNO3           ",
         "CLO             ",
         "CLOO            ",
         "CSL             ",
         "EOH             ",
         "ETHLN           ",
         "ETHN            ",
         "ETHP            ",
         "ETNO3           ",
         "ETP             ",
         "FURA            ",
         "GLYC            ",
         "GLYX            ",
         "H2O2            ",
         "HAC             ",
         "HBR             ",
         "HC5A            ",
         "HCL             ",
         "HCOOH           ",
         "HI              ",
         "HMHP            ",
         "HMML            ",
         "HNO3            ",
         "HOBR            ",
         "HOCL            ",
         "HOI             ",
         "HONIT           ",
         "HPALD1          ",
         "HPALD2          ",
         "HPALD3          ",
         "HPALD4          ",
         "HPETHNL         ",
         "I2              ",
         "I2O2            ",
         "I2O3            ",
         "I2O4            ",
         "IBR             ",
         "ICHE            ",
         "ICL             ",
         "ICN             ",
         "ICPDH           ",
         "IDC             ",
         "IDCHP           ",
         "IDHDP           ",
         "IDHPE           ",
         "IDN             ",
         "IEPOXA          ",
         "IEPOXB          ",
         "IEPOXD          ",
         "IHN1            ",
         "IHN2            ",
         "IHN3            ",
         "IHN4            ",
         "INPB            ",
         "INPD            ",
         "IONO            ",
         "IONO2           ",
         "IPRNO3          ",
         "ITCN            ",
         "ITHN            ",
         "LIMO            ",
         "LVOC            ",
         "LVOCOA          ",
         "MACR            ",
         "MACR1OOH        ",
         "MAP             ",
         "MCRDH           ",
         "MCRENOL         ",
         "MCRHN           ",
         "MCRHNB          ",
         "MCRHP           ",
         "MCT             ",
         "MEK             ",
         "MENO3           ",
         "MGLY            ",
         "MOH             ",
         "MONITS          ",
         "MONITU          ",
         "MP              ",
         "MPAN            ",
         "MPN             ",
         "MTPA            ",
         "MTPO            ",
         "MVK             ",
         "MVKDH           ",
         "MVKHC           ",
         "MVKHCB          ",
         "MVKHP           ",
         "MVKN            ",
         "MVKPC           ",
         "N2O5            ",
         "NH3             ",
         "NO2             ",
         "NPHEN           ",
         "NPRNO3          ",
         "O3              ",
         "OX              ",
         "PAN             ",
         "PHEN            ",
         "PP              ",
         "PPN             ",
         "PROPNN          ",
         "PRPN            ",
         "PRPE            ",
         "PYAC            ",
         "R4N2            ",
         "R4P             ",
         "RA3P            ",
         "RB3P            ",
         "RIPA            ",
         "RIPB            ",
         "RIPC            ",
         "RIPD            ",
         "RP              ",
         "SO2             " ;

  dfoxd = 
        1.       // ACET	      
       ,1.       // ACTA	      
       ,1.       // ALD2	      
       ,1.       // AROMP4      
       ,1.       // AROMP5      
       ,1.       // ATOOH	      
       ,1.       // BALD	      
       ,1.       // BENZP	      
       ,1.e-36   // BR2	      
       ,1.e-36   // BRCL	      
       ,1.e-36   // BRNO3	      
       ,1.       // BZCO3H      
       ,1.       // BZPAN	      
       ,1.       // CH2O	      
       ,1.e-36   // CL2	      
       ,1.e-36   // CLNO2	      
       ,1.e-36   // CLNO3	      
       ,1.e-36   // CLO	      
       ,1.e-36   // CLOO	      
       ,1.       // CSL	      
       ,1.e-36   // EOH	      
       ,1        // ETHLN	      
       ,.1       // ETHN	      
       ,.1       // ETHP	      
       ,.1       // ETNO3	      
       ,1.       // ETP
       ,1.       // FURA
       ,1.       // GLYC	      
       ,1.       // GLYX	      
       ,1.       // H2O2	      
       ,1.       // HAC	      
       ,1.e-36   // HBR	      
       ,1.e-36   // HC5A	      
       ,1.e-36   // HCL	      
       ,1.       // HCOOH	      
       ,1.e-36   // HI	      
       ,1.       // HMHP	      
       ,1.       // HMML	      
       ,1.e-36   // HNO3	      
       ,1.e-36   // HOBR	      
       ,1.e-36   // HOCL	      
       ,1.e-36   // HOI	      
       ,1.       // HONIT	      
       ,1.e-36   // HPALD1      
       ,1.e-36   // HPALD2      
       ,1.e-36   // HPALD3      
       ,1.e-36   // HPALD4      
       ,1.       // HPETHNL     
       ,1.e-36   // I2	      
       ,1.e-36   // I2O2	      
       ,1.e-36   // I2O3	      
       ,1.e-36   // I2O4	      
       ,1.e-36   // IBR	      
       ,1.       // ICHE	      
       ,1.e-36   // ICL	      
       ,1.       // ICN	      
       ,1.       // ICPDH	      
       ,1.e-36   // IDC	      
       ,1.       // IDCHP	      
       ,1.       // IDHDP	      
       ,1.       // IDHPE	      
       ,1.       // IDN	      
       ,1.       // IEPOXA      
       ,1.       // IEPOXB      
       ,1.       // IEPOXD      
       ,1.       // IHN1	      
       ,1.       // IHN2	      
       ,1.       // IHN3	      
       ,1.       // IHN4	      
       ,1.       // INPB	      
       ,1.       // INPD	      
       ,1.e-36   // IONO	      
       ,1.e-36   // IONO2	      
       ,.1       // IPRNO3      
       ,1.       // ITCN	      
       ,1.       // ITHN	      
       ,1.e-36   // LIMO	      
       ,1.       // LVOC	      
       ,1.e-36   // LVOCOA	      
       ,1        // MACR	      
       ,1        // MACR1OOH    
       ,1        // MAP	      
       ,1        // MCRDH	      
       ,1        // MCRENOL     
       ,1        // MCRHN	      
       ,1        // MCRHNB      
       ,1        // MCRHP	      
       ,1        // MCT	      
       ,1.e-36   // MEK	      
       ,.1       // MENO3	      
       ,1.       // MGLY	      
       ,1.       // MOH	      
       ,1.       // MONITS      
       ,1.       // MONITU      
       ,1.e-36   // MP	      
       ,1.       // MPAN	      
       ,1.e-36   // MPN	      
       ,1.e-36   // MTPA	      
       ,1.e-36   // MTPO	      
       ,1.       // MVK	      
       ,1.       // MVKDH	      
       ,1.       // MVKHC	      
       ,1.       // MVKHCB      
       ,1.       // MVKHP	      
       ,1.       // MVKN	      
       ,1.       // MVKPC	      
       ,1.e-36   // N2O5	      
       ,1.e-36   // NH3	      
       ,.1       // NO2	      
       ,1.       // NPHEN	      
       ,.1       // NPRNO3      
       ,1.       // O3	      
       ,1.       // OX	      
       ,1.       // PAN	      
       ,1.       // PHEN	      
       ,1.       // PP	      
       ,1.       // PPN	      
       ,1.       // PROPNN      
       ,1.e-36   // PRPE	      
       ,1.       // PRPN	      
       ,1.       // PYAC	      
       ,1.       // R4N2	      
       ,1.       // R4P	      
       ,1.       // RA3P	      
       ,1.       // RB3P	      
       ,1.       // RIPA	      
       ,1.       // RIPB	      
       ,1.       // RIPC	      
       ,1.       // RIPD	      
       ,1.       // RP	      
       ,1.e-36 ; // SO2

 dheff = 
       27.399999618530273      ,   5500.0, 0., 0., 0., 0.,  // ACET	      
       4050.0000000000000      ,   6200.0, 0., 0., 0., 0.,  // ACTA	      
       13.199999809265137      ,   5900.0, 0., 0., 0., 0.,  // ALD2	      
       410000.00000000000      ,   7500.0, 0., 0., 0., 0.,  // AROMP4      
       2000000.0000000000      ,   7500.0, 0., 0., 0., 0.,  // AROMP5      
       294.00000000000000      ,   5200.0, 0., 0., 0., 0.,  // ATOOH	      
       38.000000000000000      ,   5500.0, 0., 0., 0., 0.,  // BALD	      
       2900.0000000000000      ,   6800.0, 0., 0., 0., 0.,  // BENZP	      
      0.75999999046325684      ,   3720.0, 0., 0., 0., 0.,  // BR2	      
      0.97000002861022949      ,   5600.0, 0., 0., 0., 0.,  // BRCL	      
       0.00000000000000        ,      0.0, 0., 0., 0., 0.,  // BRNO3	      
       24000.000000000000      ,      0.0, 0., 0., 0., 0.,  // BZCO3H      
       70.000000000000000      ,   4600.0, 0., 0., 0., 0.,  // BZPAN	      
       3240.0000000000000      ,   6800.0, 0., 0., 0., 0.,  // CH2O	      
       9.2000000178813934E-002 ,   2000.0, 0., 0., 0., 0.,  // CL2	      
       0.00000000000000        ,      0.0, 0., 0., 0., 0.,  // CLNO2	      
       1.0000000200408773E+020 ,      0.0, 0., 0., 0., 0.,  // CLNO3	      
       0.00000000000000        ,      0.0, 0., 0., 0., 0.,  // CLO	      
       1.0000000000000000      ,   3500.0, 0., 0., 0., 0.,  // CLOO	      
       420.00000000000000      ,   8500.0, 0., 0., 0., 0.,  // CSL	      
       193.00000000000000      ,   6400.0, 0., 0., 0., 0.,  // EOH	      
       17000.000000000000      ,   9200.0, 0., 0., 0., 0.,  // ETHLN	      
       39000.000000000000      ,   8600.0, 0., 0., 0., 0.,  // ETHN	      
       650000.00000000000      ,   8800.0, 0., 0., 0., 0.,  // ETHP	      
       1.6000000238418579      ,   5400.0, 0., 0., 0., 0.,  // ETNO3	      
       334.00000000000000      ,   6000.0, 0., 0., 0., 0.,  // ETP	      
       1.8000000000000000E-001 ,   6100.0, 0., 0., 0., 0.,  // FURA
       41500.000000000000      ,   4600.0, 0., 0., 0., 0.,  // GLYC	      
       415000.00000000000      ,   7500.0, 0., 0., 0., 0.,  // GLYX	      
       83000.000000000000      ,   7400.0, 0., 0., 0., 0.,  // H2O2	      
       7800.0000000000000      ,      0.0, 0., 0., 0., 0.,  // HAC	      
       71000003706880.000      ,  10200.0, 0., 0., 0., 0.,  // HBR	      
       7800.0000000000000      ,      0.0, 0., 0., 0., 0.,  // HC5A	      
       62999998464.000000      ,   9000.0, 0., 0., 0., 0.,  // HCL	      
       8920.0000000000000      ,   6100.0, 0., 0., 0., 0.,  // HCOOH	      
       74299998208000.000      ,   3187.2, 0., 0., 0., 0.,  // HI	      
       1300000.0000000000      ,   5200.0, 0., 0., 0., 0.,  // HMHP	      
       120000.00000000000      ,   7200.0, 0., 0., 0., 0.,  // HMML	      
       83000.000000000000      ,   7400.0, 0., 0., 0., 0.,  // HNO3	      
       1300.0000000000000      ,   4000.0, 0., 0., 0., 0.,  // HOBR	      
       650.00000000000000      ,   5900.0, 0., 0., 0., 0.,  // HOCL	      
       15400.000000000000      ,   8371.0, 0., 0., 0., 0.,  // HOI	      
       26900000931840.000      ,   5487.0, 0., 0., 0., 0.,  // HONIT	      
       40000.000000000000      ,      0.0, 0., 0., 0., 0.,  // HPALD1      
       40000.000000000000      ,      0.0, 0., 0., 0., 0.,  // HPALD2      
       40000.000000000000      ,      0.0, 0., 0., 0., 0.,  // HPALD3      
       40000.000000000000      ,      0.0, 0., 0., 0., 0.,  // HPALD4      
       41000.000000000000      ,   4600.0, 0., 0., 0., 0.,  // HPETHNL     
       2.7000000476837158      ,   7507.4, 0., 0., 0., 0.,  // I2	      
       1.0000000200408773E+020 ,  18900.0, 0., 0., 0., 0.,  // I2O2	      
       1.0000000200408773E+020 ,  13400.0, 0., 0., 0., 0.,  // I2O3	      
       1.0000000200408773E+020 ,  13400.0, 0., 0., 0., 0.,  // I2O4	      
       24.000000000000000      ,   4916.7, 0., 0., 0., 0.,  // IBR	      
       80000000.000000000      ,      0.0, 0., 0., 0., 0.,  // ICHE	      
       111.00000000000000      ,   2105.5, 0., 0., 0., 0.,  // ICL	      
       17000.000000000000      ,   9200.0, 0., 0., 0., 0.,  // ICN	      
       100000000.00000000      ,   7200.0, 0., 0., 0., 0.,  // ICPDH	      
       40000.000000000000      ,      0.0, 0., 0., 0., 0.,  // IDC	      
       100000000.00000000      ,   7200.0, 0., 0., 0., 0.,  // IDCHP	      
       100000000.00000000      ,   7200.0, 0., 0., 0., 0.,  // IDHDP	      
       100000000.00000000      ,   7200.0, 0., 0., 0., 0.,  // IDHPE	      
       100000000.00000000      ,   7200.0, 0., 0., 0., 0.,  // IDN	      
       80000000.000000000      ,      0.0, 0., 0., 0., 0.,  // IEPOXA      
       80000000.000000000      ,      0.0, 0., 0., 0., 0.,  // IEPOXB      
       80000000.000000000      ,      0.0, 0., 0., 0., 0.,  // IEPOXD      
       17000.000000000000      ,   9200.0, 0., 0., 0., 0.,  // IHN1	      
       17000.000000000000      ,   9200.0, 0., 0., 0., 0.,  // IHN2	      
       17000.000000000000      ,   9200.0, 0., 0., 0., 0.,  // IHN3	      
       17000.000000000000      ,   9200.0, 0., 0., 0., 0.,  // IHN4	      
       17000.000000000000      ,   9200.0, 0., 0., 0., 0.,  // INPB	      
       17000.000000000000      ,   9200.0, 0., 0., 0., 0.,  // INPD	      
      0.30000001192092896      ,   7240.4, 0., 0., 0., 0.,  // IONO	      
       1.0000000200408773E+020 ,   3980.0, 0., 0., 0., 0.,  // IONO2	      
      0.79000002145767212      ,   5400.0, 0., 0., 0., 0.,  // IPRNO3      
       100000000.00000000      ,   7200.0, 0., 0., 0., 0.,  // ITCN	      
       100000000.00000000      ,   7200.0, 0., 0., 0., 0.,  // ITHN	      
       7.0000000298023224E-002 ,      0.0, 0., 0., 0., 0.,  // LIMO	      
       100000000.00000000      ,   7200.0, 0., 0., 0., 0.,  // LVOC	      
       0.00000000000000        ,      0.0, 0., 0., 0., 0.,  // LVOCOA	      
       4.8600001335144043      ,   4300.0, 0., 0., 0., 0.,  // MACR	      
       294.00000000000000      ,   5200.0, 0., 0., 0., 0.,  // MACR1OOH    
       840.00000000000000      ,   5300.0, 0., 0., 0., 0.,  // MAP	      
       1400000.0000000000      ,   7200.0, 0., 0., 0., 0.,  // MCRDH	      
       294.00000000000000      ,   5200.0, 0., 0., 0., 0.,  // MCRENOL     
       17000.000000000000      ,   9200.0, 0., 0., 0., 0.,  // MCRHN	      
       17000.000000000000      ,   9200.0, 0., 0., 0., 0.,  // MCRHNB      
       1400000.0000000000      ,   7200.0, 0., 0., 0., 0.,  // MCRHP	      
       420.00000000000000      ,   8500.0, 0., 0., 0., 0.,  // MCT	      
       18.200000000000000      ,   5700.0, 0., 0., 0., 0.,  // MEK	      
       11.000000000000000      ,   4700.0, 0., 0., 0., 0.,  // MENO3	      
       32400.000000000000      ,   6200.0, 0., 0., 0., 0.,  // MGLY	      
       203.00000000000000      ,   5600.0, 0., 0., 0., 0.,  // MOH	      
       17000.000000000000      ,   9200.0, 0., 0., 0., 0.,  // MONITS      
       17000.000000000000      ,   9200.0, 0., 0., 0., 0.,  // MONITU      
       294.00000000000000      ,   5200.0, 0., 0., 0., 0.,  // MP	      
       1.7200000286102295      ,      0.0, 0., 0., 0., 0.,  // MPAN	      
       294.00000000000000      ,   5200.0, 0., 0., 0., 0.,  // MPN	      
       4.8999998718500137E-002 ,      0.0, 0., 0., 0., 0.,  // MTPA	      
       4.8999998718500137E-002 ,      0.0, 0., 0., 0., 0.,  // MTPO	      
       26.299999237060547      ,   4800.0, 0., 0., 0., 0.,  // MVK	      
       1400000.0000000000      ,   7200.0, 0., 0., 0., 0.,  // MVKDH	      
       1400000.0000000000      ,   7200.0, 0., 0., 0., 0.,  // MVKHC	      
       1400000.0000000000      ,   7200.0, 0., 0., 0., 0.,  // MVKHCB      
       1400000.0000000000      ,   7200.0, 0., 0., 0., 0.,  // MVKHP	      
       17000.000000000000      ,   9200.0, 0., 0., 0., 0.,  // MVKN	      
       1400000.0000000000      ,   7200.0, 0., 0., 0., 0.,  // MVKPC	      
       0.0000000000000000      ,      0.0, 0., 0., 0., 0.,  // N2O5	      
       3300000.0000000000      ,   4100.0, 0., 0., 0., 0.,  // NH3	      
       0.0000000000000000      ,      0.0, 0., 0., 0., 0.,  // NO2	      
       2300.0000000000000      ,      0.0, 0., 0., 0., 0.,  // NPHEN	      
       1.1000000238418579      ,   5500.0, 0., 0., 0., 0.,  // NPRNO3      
       1.0132499970495701E-002 ,   2800.0, 0., 0., 0., 0.,  // O3	      
       1.0132499970495701E-002 ,   2800.0, 0., 0., 0., 0.,  // OX	      
       2.940000572204590       ,   5700.0, 0., 0., 0., 0.,  // PAN	      
       2800.0000000000000      ,   2700.0, 0., 0., 0., 0.,  // PHEN	      
       294.00000000000000      ,   5200.0, 0., 0., 0., 0.,  // PP	      
       2.9400000572204590      ,      0.0, 0., 0., 0., 0.,  // PPN	      
       1000.0000000000000      ,      0.0, 0., 0., 0., 0.,  // PROPNN      
       7.4000000000000000E-003 ,   3400.0, 0., 0., 0., 0.,  // PRPE	      
       294.00000000000000      ,   5200.0, 0., 0., 0., 0.,  // PRPN	      
       314000.00000000000      ,   5100.0, 0., 0., 0., 0.,  // PYAC	      
       1.0000000000000000      ,   5800.0, 0., 0., 0., 0.,  // R4N2	      
       294.00000000000000      ,   5200.0, 0., 0., 0., 0.,  // R4P	      
       294.00000000000000      ,   5200.0, 0., 0., 0., 0.,  // RA3P	      
       294.00000000000000      ,   5200.0, 0., 0., 0., 0.,  // RB3P	      
       1700000.0000000000      ,      0.0, 0., 0., 0., 0.,  // RIPA	      
       1700000.0000000000      ,      0.0, 0., 0., 0., 0.,  // RIPB	      
       1700000.0000000000      ,      0.0, 0., 0., 0., 0.,  // RIPC	      
       1700000.0000000000      ,      0.0, 0., 0., 0., 0.,  // RIPD	      
       294.00000000000000      ,   5200.0, 0., 0., 0., 0.,  // RP	      
       0.0000000000000000      ,      0.0, 0., 0., 0., 0. ; // SO2         

  mol_wghts =
         ,58.090000000000003   // ACET	      
         ,60.060000000000002   // ACTA	      
         ,44.060000000000002   // ALD2	      
         ,68.079999999999998   // AROMP4      
         ,98.099999999999994   // AROMP5      
         ,90.090000000000003   // ATOOH	      
         ,106.12000000000000   // BALD	      
         ,110.11000000000000   // BENZP	      
         ,159.80000000000001   // BR2	      
         ,115.45000000000000   // BRCL	      
         ,141.91000000000000   // BRNO3	      
         ,138.12000000000000   // BZCO3H      
         ,183.12000000000000   // BZPAN	      
         ,30.030000000000001   // CH2O	      
         ,70.900000000000006   // CL2	      
         ,81.450000000000003   // CLNO2	      
         ,97.450000000000003   // CLNO3	      
         ,51.450000000000003   // CLO	      
         ,67.450000000000003   // CLOO	      
         ,108.14000000000000   // CSL	      
         ,46.070000000000000   // EOH	      
         ,105.06000000000000   // ETHLN	      
         ,107.06999999999999   // ETHN	      
         ,78.069999999999993   // ETHP	      
         ,91.079999999999998   // ETNO3	      
         ,62.079999999999998   // ETP	      
         ,68.070000000000000   // FURA
	 ,60.060000000000002   // GLYC	      
         ,58.039999999999999   // GLYX	      
         ,34.020000000000003   // H2O2	      
         ,74.079999999999998   // HAC	      
         ,80.909999999999997   // HBR	      
         ,100.13000000000000   // HC5A	      
         ,36.450000000000003   // HCL	      
         ,46.030000000000001   // HCOOH	      
         ,127.91000000000000   // HI	      
         ,64.049999999999997   // HMHP	      
         ,102.09999999999999   // HMML	      
         ,63.009999999999998   // HNO3	      
         ,96.909999999999997   // HOBR	      
         ,52.450000000000003   // HOCL	      
         ,143.88999999999999   // HOI	      
         ,215.00000000000000   // HONIT	      
         ,116.13000000000000   // HPALD1      
         ,116.13000000000000   // HPALD2      
         ,116.13000000000000   // HPALD3      
         ,116.13000000000000   // HPALD4      
         ,76.060000000000002   // HPETHNL     
         ,253.80000000000001   // I2	      
         ,285.80000000000001   // I2O2	      
         ,301.80000000000001   // I2O3	      
         ,317.80000000000001   // I2O4	      
         ,206.90000000000001   // IBR	      
         ,116.13000000000000   // ICHE	      
         ,162.44999999999999   // ICL	      
         ,145.13000000000000   // ICN	      
         ,150.15000000000001   // ICPDH	      
         ,98.109999999999999   // IDC	      
         ,148.13000000000000   // IDCHP	      
         ,168.16999999999999   // IDHDP	      
         ,150.15000000000001   // IDHPE	      
         ,192.15000000000001   // IDN	      
         ,106.14000000000000   // IEPOXA      
         ,106.14000000000000   // IEPOXB      
         ,106.14000000000000   // IEPOXD      
         ,147.15000000000001   // IHN1	      
         ,147.15000000000001   // IHN2	      
         ,147.15000000000001   // IHN3	      
         ,147.15000000000001   // IHN4	      
         ,163.15000000000001   // INPB	      
         ,163.15000000000001   // INPD	      
         ,172.91000000000000   // IONO	      
         ,188.91000000000000   // IONO2	      
         ,105.11000000000000   // IPRNO3      
         ,195.15000000000000   // ITCN	      
         ,197.16999999999999   // ITHN	      
         ,136.25999999999999   // LIMO	      
         ,154.19000000000000   // LVOC	      
         ,154.19000000000000   // LVOCOA
         ,70.099999999999994   // MACR	      
         ,102.09999999999999   // MACR1OOH    
         ,76.060000000000002   // MAP	      
         ,104.12000000000000   // MCRDH	      
         ,86.099999999999994   // MCRENOL     
         ,149.11000000000001   // MCRHN	      
         ,149.11000000000001   // MCRHNB      
         ,120.12000000000000   // MCRHP	      
         ,124.00000000000000   // MCT	      
         ,72.110000000000000   // MEK	      
         ,77.049999999999997   // MENO3	      
         ,72.069999999999993   // MGLY	      
         ,32.049999999999997   // MOH	      
         ,215.28000000000000   // MONITS      
         ,215.28000000000000   // MONITU      
         ,48.050000000000000   // MP	      
         ,147.09999999999999   // MPAN	      
         ,93.050000000000000   // MPN	      
         ,136.25999999999999   // MTPA	      
         ,136.25999999999999   // MTPO	      
         ,70.090000000000003   // MVK	      
         ,105.13000000000000   // MVKDH	      
         ,102.09999999999999   // MVKHC	      
         ,102.09999999999999   // MVKHCB      
         ,120.12000000000000   // MVKHP	      
         ,149.12000000000000   // MVKN	      
         ,118.09999999999999   // MVKPC	      
         ,108.02000000000000   // N2O5	      
         ,17.039999999999999   // NH3	      
         ,46.009999999999998   // NO2	      
         ,139.11000000000001   // NPHEN	      
         ,105.11000000000000   // NPRNO3      
         ,48.000000000000000   // O3	      
         ,48.000000000000000   // OX	      
         ,121.06000000000000   // PAN	      
         ,94.109999999999999   // PHEN	      
         ,92.109999999999999   // PP	      
         ,135.08000000000001   // PPN	      
         ,119.08000000000000   // PROPNN      
         ,42.090000000000000   // PRPE	      
         ,137.11000000000001   // PRPN	      
         ,88.069999999999993   // PYAC	      
         ,119.09999999999999   // R4N2	      
         ,90.140000000000001   // R4P	      
         ,76.109999999999999   // RA3P	      
         ,76.109999999999999   // RB3P	      
         ,118.15000000000001   // RIPA	      
         ,118.15000000000001   // RIPB	      
         ,118.15000000000001   // RIPC	      
         ,118.15000000000001   // RIPD	      
         ,90.090000000000003   // RP	      
         ,64.040000000000006 ; // SO2         

}